library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


Entity VGA_tb is
end VGA_tb;

Architecture behavioral of VGA_tb is
begin

end behavioral;
